module stickman (
    input  wire [6:0] y,       // Row index (0–15)
    output wire [127:0] row     // 16-bit row data
);

    reg [127:0] sprite_rom [0:127];

    initial begin
    sprite_rom[0] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 0
    sprite_rom[1] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 1
    sprite_rom[2] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 2
    sprite_rom[3] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 3
    sprite_rom[4] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 4
    sprite_rom[5] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 5
    sprite_rom[6] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 6
    sprite_rom[7] = 128'b00000000000000000000000000111111111111111000000000000000000000000000000000000001111111111111100000000000000000000000000000000000;  // row 7
    sprite_rom[8] = 128'b00000000000000000000000000111111111111111000000000000000000000000000000000000001111111111111100000000000000000000000000000000000;  // row 8
    sprite_rom[9] = 128'b00000000000000000000000000111111111111111000000000000000000000000000000000000001111111111111100000000000000000000000000000000000;  // row 9
    sprite_rom[10] = 128'b00000000000000000000000000111111111111111000000000000000000000000000000000000001111111111111100000000000000000000000000000000000;  // row 10
    sprite_rom[11] = 128'b00000000000000000000001111111111111111111000011111111111111111111111111111111111111111111111111110000000000000000000000000000000;  // row 11
    sprite_rom[12] = 128'b00000000000000000000001111111111111111111000011111111111111111111111111111111111111111111111111110000000000000000000000000000000;  // row 12
    sprite_rom[13] = 128'b00000000000000000000001111111111111111111000011111111111111111111111111111111111111111111111111110000000000000000000000000000000;  // row 13
    sprite_rom[14] = 128'b00000000000000000000001111111111111111111000011111111111111111111111111111111111111111111111111110000000000000000000000000000000;  // row 14
    sprite_rom[15] = 128'b00000000000000000000001111111111111111111111100000000000000000000000000000011111111111111111111110000000000000000000000000000000;  // row 15
    sprite_rom[16] = 128'b00000000000000000000001111111111111111111111100000000000000000000000000000011111111111111111111110000000000000000000000000000000;  // row 16
    sprite_rom[17] = 128'b00000000000000000000001111111111111111111111100000000000000000000000000000011111111111111111111110000000000000000000000000000000;  // row 17
    sprite_rom[18] = 128'b00000000000000000000001111111111111111111111100000000000000000000000000000011111111111111111111110000000000000000000000000000000;  // row 18
    sprite_rom[19] = 128'b00000000000000000000001111111111111111111000000000000000000000000000000000000000000111111111111110000000000000000000000000000000;  // row 19
    sprite_rom[20] = 128'b00000000000000000000001111111111111111111000000000000000000000000000000000000000000111111111111110000000000000000000000000000000;  // row 20
    sprite_rom[21] = 128'b00000000000000000000001111111111111111111000000000000000000000000000000000000000000111111111111110000000000000000000000000000000;  // row 21
    sprite_rom[22] = 128'b00000000000000000000001111111111111111111000000000000000000000000000000000000000000111111111111110000000000000000000000000000000;  // row 22
    sprite_rom[23] = 128'b00000000000000000000001111111111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000;  // row 23
    sprite_rom[24] = 128'b00000000000000000000001111111111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000;  // row 24
    sprite_rom[25] = 128'b00000000000000000000001111111111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000;  // row 25
    sprite_rom[26] = 128'b00000000000000000000001111111111111110000000000000000000000000000000000000000000000000000111111110000000000000000000000000000000;  // row 26
    sprite_rom[27] = 128'b00000000000000000000000000111111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000;  // row 27
    sprite_rom[28] = 128'b00000000000000000000000000111111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000;  // row 28
    sprite_rom[29] = 128'b00000000000000000000000000111111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000;  // row 29
    sprite_rom[30] = 128'b00000000000000000000000000111111100000000000000000000000000000000000000000000000000000000111100000000000000000000000000000000000;  // row 30
    sprite_rom[31] = 128'b00000000000000000000001111111000000000000000011111111111100000000000000000000000000000111111100000000000000000000000000000000000;  // row 31
    sprite_rom[32] = 128'b00000000000000000000001111111000000000000000011111111111100000000000000000000000000000111111100000000000000000000000000000000000;  // row 32
    sprite_rom[33] = 128'b00000000000000000000001111111000000000000000011111111111100000000000000000000000000000111111100000000000000000000000000000000000;  // row 33
    sprite_rom[34] = 128'b00000000000000000000001111111000000000000000011111111111100000000000000000000000000000111111100000000000000000000000000000000000;  // row 34
    sprite_rom[35] = 128'b00000000000000000000001111111000000000000111111111111111111110000000000000000000000111111111100000000000000000000000000000000000;  // row 35
    sprite_rom[36] = 128'b00000000000000000000001111111000000000000111111111111111111110000000000000000000000111111111100000000000000000000000000000000000;  // row 36
    sprite_rom[37] = 128'b00000000000000000000001111111000000000000111111111111111111110000000000000000000000111111111100000000000000000000000000000000000;  // row 37
    sprite_rom[38] = 128'b00000000000000000000001111111000000000000111111111111111111110000000000000000000000111111111100000000000000000000000000000000000;  // row 38
    sprite_rom[39] = 128'b00000000000000000000001111111000000000000111111111111000011111111000000000000001111111000111100000000000000000000000000000000000;  // row 39
    sprite_rom[40] = 128'b00000000000000000000001111111000000000000111111111111000011111111000000000000001111111000111100000000000000000000000000000000000;  // row 40
    sprite_rom[41] = 128'b00000000000000000000001111111000000000000111111111111000011111111000000000000001111110000111100000000000000000000000000000000000;  // row 41
    sprite_rom[42] = 128'b00000000000000000000001111111000000000000111111111111000011111111000000000000001111110000111100000000000000000000000000000000000;  // row 42
    sprite_rom[43] = 128'b00000000000000000000001111111000000000000111111111111000011111111000000000000001111110000111100000000000000000000000000000000000;  // row 43
    sprite_rom[44] = 128'b00000000000000000000001111111000000000000111111111111000011111111000000000000001111110000111100000000000000000000000000000000000;  // row 44
    sprite_rom[45] = 128'b00000000000000000000001111111000000000000111111111111000011111111000000000000001111110000111100000000000000000000000000000000000;  // row 45
    sprite_rom[46] = 128'b00000000000000000000001111111000000000000111111111111000011111111000000000000001111110000111100000000000000000000000000000000000;  // row 46
    sprite_rom[47] = 128'b00000000000000000000001111111000000000000000011111111111111110000000000000000000000111111111100000000000000000000000000000000000;  // row 47
    sprite_rom[48] = 128'b00000000000000000000001111111000000000000000011111111111111110000000000000000000000111111111100000000000000000000000000000000000;  // row 48
    sprite_rom[49] = 128'b00000000000000000000001111111000000000000000011111111111111110000000000000000000000111111111100000000000000000000000000000000000;  // row 49
    sprite_rom[50] = 128'b00000000000000000000001111111000000000000000011111111111111110000000000000000000000111111111100000000000000000000000000000000000;  // row 50
    sprite_rom[51] = 128'b00000000000000000000001111111000000000000000000000000000000000000000000111111111111000000111100000000000000000000000000000000000;  // row 51
    sprite_rom[52] = 128'b00000000000000000000001111111000000000000000000000000000000000000000000111111111111000000111100000000000000000000000000000000000;  // row 52
    sprite_rom[53] = 128'b00000000000000000000001111111000000000000000000000000000000000000000000111111111111000000111100000000000000000000000000000000000;  // row 53
    sprite_rom[54] = 128'b00000000000000000000001111111000000000000000000000000000000000000000000111111111111000000111100000000000000000000000000000000000;  // row 54
    sprite_rom[55] = 128'b00000000000000000000000000111111100000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000;  // row 55
    sprite_rom[56] = 128'b00000000000000000000000000111111100000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000;  // row 56
    sprite_rom[57] = 128'b00000000000000000000000000111111100000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000;  // row 57
    sprite_rom[58] = 128'b00000000000000000000000000111111100000000000000000000000000000000000000000011110000000000111100000000000000000000000000000000000;  // row 58
    sprite_rom[59] = 128'b00000000000000000000000000000111111111111000000000000000000000011111111111111110000000111000000000000000000000000000000000000000;  // row 59
    sprite_rom[60] = 128'b00000000000000000000000000000111111111111000000000000000000000011111111111111110000000111000000000000000000000000000000000000000;  // row 60
    sprite_rom[61] = 128'b00000000000000000000000000000111111111111000000000000000000000011111111111111110000000111000000000000000000000000000000000000000;  // row 61
    sprite_rom[62] = 128'b00000000000000000000000000000111111111111000000000000000000000011111111111111110000000111000000000000000000000000000000000000000;  // row 62
    sprite_rom[63] = 128'b00000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000;  // row 63
    sprite_rom[64] = 128'b00000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000;  // row 64
    sprite_rom[65] = 128'b00000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000;  // row 65
    sprite_rom[66] = 128'b00000000000000000000000000111111111111111111111110000000000000000000000000000001111111111111111111100000000000000000000000000000;  // row 66
    sprite_rom[67] = 128'b00000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000;  // row 67
    sprite_rom[68] = 128'b00000000000000000000001111111111111111111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000;  // row 68
    sprite_rom[69] = 128'b00000000000000000000001111111111111111111111111111111111111111111111111111111111111111100001111111111110000000000000000000000000;  // row 69
    sprite_rom[70] = 128'b00000000000000000000001111111111111111111111111111111111111111111111111111111111111111100001111111111110000000000000000000000000;  // row 70
    sprite_rom[71] = 128'b00000000000000000011111111111111111111111111111111111111111111111111111111111111111111100111111111111110000000000000000000000000;  // row 71
    sprite_rom[72] = 128'b00000000000000000011111111111111111111111111111111111111111111111111111111111111111111100111111111111110000000000000000000000000;  // row 72
    sprite_rom[73] = 128'b00000000000000000011111111111111111111111111111111111111111111111111111111111111111111100111111111111110000000000000000000000000;  // row 73
    sprite_rom[74] = 128'b00000000000000000011111111111111111111111111111111111111111111111111111111111111111111100111111111111110000000000000000000000000;  // row 74
    sprite_rom[75] = 128'b00000000000000000011111111111111111110000111111111111000000000000000000000000001111111100111111111111110000000000000000000000000;  // row 75
    sprite_rom[76] = 128'b00000000000000000011111111111111111110000111111111111000000000000000000000000001111111100111111111111110000000000000000000000000;  // row 76
    sprite_rom[77] = 128'b00000000000000000011111111111111111110000111111111111000000000000000000000000001111111100111111111111110000000000000000000000000;  // row 77
    sprite_rom[78] = 128'b00000000000000000011111111111111111110000111111111111000000000000000000000000001111111100111111111111110000000000000000000000000;  // row 78
    sprite_rom[79] = 128'b00000000000000000011111111111111100001111111100000000000000000000000000000000000000111111111111111111110000000000000000000000000;  // row 79
    sprite_rom[80] = 128'b00000000000000000011111111111111100001111111100000000000000000000000000000000000000111111111111111111110000000000000000000000000;  // row 80
    sprite_rom[81] = 128'b00000000000000000011111111111111100001111111100000000000000000000000000000000000000111111111111111111110000000000000000000000000;  // row 81
    sprite_rom[82] = 128'b00000000000000000011111111111111100001111111100000000000000000000000000000000000000111111111111111111110000000000000000000000000;  // row 82
    sprite_rom[83] = 128'b00000000000000000011111111111111111111111000000000000000000000000000000000000000000111111111111111100000000000000000000000000000;  // row 83
    sprite_rom[84] = 128'b00000000000000000011111111111111111111111000000000000000000000000000000000000000000111111111111111100000000000000000000000000000;  // row 84
    sprite_rom[85] = 128'b00000000000000000011111111111111111111111000000000000000000000000000000000000000000111111111111111100000000000000000000000000000;  // row 85
    sprite_rom[86] = 128'b00000000000000000011111111111111111111111000000000000000000000000000000000000000000111111111111111100000000000000000000000000000;  // row 86
    sprite_rom[87] = 128'b00000000000000000000001111111111111111111000000000000000000000000000000000000000000111100000000000000000000000000000000000000000;  // row 87
    sprite_rom[88] = 128'b00000000000000000000001111111111111111111000000000000000000000000000000000000000000111100000000000000000000000000000000000000000;  // row 88
    sprite_rom[89] = 128'b00000000000000000000001111111111111111111000000000000000000000000000000000000000000111100000000000000000000000000000000000000000;  // row 89
    sprite_rom[90] = 128'b00000000000000000000001111111111111111111000000000000000000000000000000000000000000111100000000000000000000000000000000000000000;  // row 90
    sprite_rom[91] = 128'b00000000000000000000000000111111111110000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000;  // row 91
    sprite_rom[92] = 128'b00000000000000000000000000111111111110000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000;  // row 92
    sprite_rom[93] = 128'b00000000000000000000000000111111111110000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000;  // row 93
    sprite_rom[94] = 128'b00000000000000000000000000111111111110000000000000000000000000000000000000000000000111100000000000000000000000000000000000000000;  // row 94
    sprite_rom[95] = 128'b00000000000000000000000000000111111111111000000000000000000000000000000000000001111111111110000000000000000000000000000000000000;  // row 95
    sprite_rom[96] = 128'b00000000000000000000000000000111111111111000000000000000000000000000000000000001111111111110000000000000000000000000000000000000;  // row 96
    sprite_rom[97] = 128'b00000000000000000000000000000111111111111000000000000000000000000000000000000001111111111110000000000000000000000000000000000000;  // row 97
    sprite_rom[98] = 128'b00000000000000000000000000000111111111111000000000000000000000000000000000000001111111111110000000000000000000000000000000000000;  // row 98
    sprite_rom[99] = 128'b00000000000000000000000000000111111111111111100000000000000000000000000000011111111111111110000000000000000000000000000000000000;  // row 99
    sprite_rom[100] = 128'b00000000000000000000000000000111111111111111100000000000000000000000000000011111111111111110000000000000000000000000000000000000;  // row 100
    sprite_rom[101] = 128'b00000000000000000000000000000111111111111111100000000000000000000000000000011111111111111110000000000000000000000000000000000000;  // row 101
    sprite_rom[102] = 128'b00000000000000000000000000000111111111111111100000000000000000000000000000011111111111111110000000000000000000000000000000000000;  // row 102
    sprite_rom[103] = 128'b00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000;  // row 103
    sprite_rom[104] = 128'b00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000;  // row 104
    sprite_rom[105] = 128'b00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000;  // row 105
    sprite_rom[106] = 128'b00000000000000000000000001111111111111111111111111111111111111111111111111111111111111111110000000000000000000000000000000000000;  // row 106
    sprite_rom[107] = 128'b00000000000000000000000001111111111111111111111111111000000000000001111111111111111111111110000000000000000000000000000000000000;  // row 107
    sprite_rom[108] = 128'b00000000000000000000000001111111111111111111111111111000000000000001111111111111111111111110000000000000000000000000000000000000;  // row 108
    sprite_rom[109] = 128'b00000000000000000000000001111111111111111111111111111000000000000001111111111111111111111110000000000000000000000000000000000000;  // row 109
    sprite_rom[110] = 128'b00000000000000000000000001111111111111111111111111111000000000000001111111111111111111111110000000000000000000000000000000000000;  // row 110
    sprite_rom[111] = 128'b00000000000000000000000001111111111111111111100000000000000000000000000111111111111111111111111000000000000000000000000000000000;  // row 111
    sprite_rom[112] = 128'b00000000000000000000000001111111111111111111100000000000000000000000000111111111111111111111111000000000000000000000000000000000;  // row 112
    sprite_rom[113] = 128'b00000000000000000000000001111111111111111111100000000000000000000000000111111111111111111111111000000000000000000000000000000000;  // row 113
    sprite_rom[114] = 128'b00000000000000000000000001111111111111111111100000000000000000000000000111111111111111111111111000000000000000000000000000000000;  // row 114
    sprite_rom[115] = 128'b00000000000000000000000001111111111111111000000000000000000000000000000111111111111111111111111111100000000000000000000000000000;  // row 115
    sprite_rom[116] = 128'b00000000000000000000000001111111111111111000000000000000000000000000000111111111111111111111111111100000000000000000000000000000;  // row 116
    sprite_rom[117] = 128'b00000000000000000000000001111111111111111000000000000000000000000000000111111111111111111111111111100000000000000000000000000000;  // row 117
    sprite_rom[118] = 128'b00000000000000000000000001111111111111111000000000000000000000000000000111111111111111111111111111100000000000000000000000000000;  // row 118
    sprite_rom[119] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 119
    sprite_rom[120] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 120
    sprite_rom[121] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 121
    sprite_rom[122] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 122
    sprite_rom[123] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 123
    sprite_rom[124] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 124
    sprite_rom[125] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 125
    sprite_rom[126] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 126
    sprite_rom[127] = 128'b00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;  // row 127
    end

    assign row = sprite_rom[y];

endmodule
